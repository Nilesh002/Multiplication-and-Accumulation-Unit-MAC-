module adder24(a,b,s);
input [23:0]a,b;
output [23:0]s;

assign s=a+b;

endmodule
