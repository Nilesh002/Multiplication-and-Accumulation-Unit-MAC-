module add48(a,b,s);
input [47:0]a,b;
output [47:0]s;

assign s=a+b;

endmodule
